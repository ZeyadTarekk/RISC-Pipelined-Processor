module IdExBuffer (
    input RegWrite,
    MemOrReg,
    DestOrPrivate,
    MemWrite,
    MemRead,
    clk,
    SPOrALUres,
    immOrReg,
    updateStatus,
    BranchFlag,
		makeMeBubble,

    input [3:0] regDestAddress, regSrcAddress, AlUControl,
    input [2:0] funCode,
    input [15:0] RegSrc, RegDest, imm,
    input [1:0] SPOpeartion, carryFlag,
		
    output reg oRegWrite,
    oMemOrReg,
    oMemWrite,
    oMemRead,
    oDestOrPrivate,
    oSPOrALUres,
    oimmOrReg,
    oupdateStatus,
    oBranchFlag,
    output reg [3:0] oRegDestAddress, oRegSrcAddress, oAlUControl,
    output reg [15:0] oRegSrc, oRegDest, oimm,
    output reg [1:0] oSPOpeartion, ocarryFlag,
    output reg [2:0] ofunCode
);

  initial begin
    oRegWrite = 0;
    oMemOrReg = 0;
    oDestOrPrivate = 0;
    oRegDestAddress = 0;
    oRegSrcAddress = 0;
    oSPOpeartion = 0;
    oMemWrite = 0;
    oMemRead = 0;
    oSPOrALUres = 0;
    oRegSrc = 0;
    oRegDest = 0;
    oimmOrReg = 0;
    oupdateStatus = 0;
    oAlUControl = 0;
    ocarryFlag = 0;
    ofunCode = 0;
    oimm = 0;
    oBranchFlag = 0;
  end

  always @(posedge clk) begin
    oRegWrite = RegWrite;
    oMemOrReg = MemOrReg;
    oDestOrPrivate = DestOrPrivate;
    oSPOpeartion = SPOpeartion;
    oMemWrite = MemWrite;
    oMemRead = MemRead;
    oSPOrALUres = SPOrALUres;
    oRegSrc = RegSrc;
    oRegDest = RegDest;
    oimmOrReg = immOrReg;
    oupdateStatus = updateStatus;
    oAlUControl = AlUControl;
    ocarryFlag = carryFlag;
    ofunCode = funCode;
    oimm = imm;
    oBranchFlag = BranchFlag;

		if (makeMeBubble == 1'b1) begin
			oRegDestAddress = 4'b1111;
			oRegSrcAddress = 4'b1111;
		end else begin
			oRegDestAddress = regDestAddress;
			oRegSrcAddress = regSrcAddress;
		end
  end

endmodule
